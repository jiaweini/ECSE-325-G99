library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use STD.textio.all;
use ieee.std_logic_textio.all;

entit g99_MAC_tb is
end g99_MAC_tb;

architecture test of g99_MAC_tb is
component g99_MAC is
port (x		: in	std_logic_vector(down to);



)




begin
end architecture test;